--* ><(((('> * Puli puli * ><(((('> // Ƹ̵̡Ӝ̵̨̄Ʒ * swish swish* Ƹ̵̡Ӝ̵̨̄Ʒ Ƹ̵̡Ӝ̵̨̄Ʒ // (っ◕‿◕)╭∩╮^H^H^Hっ
LIBRARY ieee;USE ieee.std_logic_1164.all;USE ieee.std_logic_arith.all;ENTITY reg_bank_1col IS PORT(clk:IN std_logic;nullify:IN std_logic;pixd_in:IN std_logic_vector(23 DOWNTO 0);rst_n:IN std_logic;write:IN std_logic;y:IN std_logic_vector(7 DOWNTO 0);pixd_out:OUT std_logic_vector(23 DOWNTO 0));END reg_bank_1col ;LIBRARY ieee;USE ieee.std_logic_1164.all;USE ieee.std_logic_arith.all;ARCHITECTURE struct OF reg_bank_1col IS SIGNAL z60a67f27d:std_logic_vector(23 DOWNTO 0);SIGNAL zc44f0ab3b:std_logic_vector(23 DOWNTO 0);SIGNAL ze64054cb6:std_logic_vector(23 DOWNTO 0);SIGNAL z508ec0017:std_logic;SIGNAL z1934d98a3:std_logic;SIGNAL zb48298c48:std_logic;SIGNAL z9f041aaff:std_logic;SIGNAL zcf058ee7c:std_logic;SIGNAL ze6d31b4ac:std_logic;SIGNAL z1b791bfd5:std_logic;SIGNAL z45a1dff88:std_logic;SIGNAL zc83e54d35:std_logic;SIGNAL z22f92b4dd:std_logic_vector(3 DOWNTO 0);SIGNAL z197a0495d:std_logic_vector(2 DOWNTO 0);SIGNAL z75dc1577a:std_logic;SIGNAL z833ab3bd5:std_logic;SIGNAL zc57c46db4:std_logic;SIGNAL z1ea89dc0d:std_logic;SIGNAL zcd48e1f4f:std_logic;SIGNAL z36424fa31:std_logic;SIGNAL z0068e7d64:std_logic;SIGNAL zb30429bb4:std_logic;SIGNAL z564ee05a3:std_logic_vector(23 DOWNTO 0);SIGNAL z0a9315da3:std_logic_vector(23 DOWNTO 0);SIGNAL z6bb6c7052:std_logic_vector(23 DOWNTO 0);SIGNAL z163c5325c:std_logic_vector(23 DOWNTO 0);SIGNAL z84b2eb77e:std_logic_vector(23 DOWNTO 0);SIGNAL zf5226fb5c:std_logic_vector(7 DOWNTO 0);COMPONENT reg_bank_1px PORT(clk:IN std_logic ;nullify:IN std_logic ;pixd_in:IN std_logic_vector(23 DOWNTO 0);rst_n:IN std_logic ;write:IN std_logic ;pixd_out:OUT std_logic_vector(23 DOWNTO 0));END COMPONENT;BEGIN zc57c46db4<=write AND z1934d98a3;z1ea89dc0d<=write AND zb48298c48;zcd48e1f4f<=write AND z75dc1577a;z36424fa31<=write AND z833ab3bd5;z508ec0017<=write AND z0068e7d64;ze6d31b4ac<=write AND zb30429bb4;z1b791bfd5<=write AND z9f041aaff;z45a1dff88<=write AND zcf058ee7c;zc83e54d35<='1';zf57631b0a:PROCESS(zc83e54d35, y)BEGIN IF(y(0)=zc83e54d35)THEN z22f92b4dd<="0000";ELSIF(y(1)=zc83e54d35)THEN z22f92b4dd<="0001";ELSIF(y(2)=zc83e54d35)THEN z22f92b4dd<="0010";ELSIF(y(3)=zc83e54d35)THEN z22f92b4dd<="0011";ELSIF(y(4)=zc83e54d35)THEN z22f92b4dd<="0100";ELSIF(y(5)=zc83e54d35)THEN z22f92b4dd<="0101";ELSIF(y(6)=zc83e54d35)THEN z22f92b4dd<="0110";ELSIF(y(7)=zc83e54d35)THEN z22f92b4dd<="0111";ELSE z22f92b4dd<="1000";END IF;END PROCESS zf57631b0a;z197a0495d<=z22f92b4dd(2)& z22f92b4dd(1)& z22f92b4dd(0);z7d086e91c:PROCESS(z163c5325c, z6bb6c7052, z0a9315da3, z564ee05a3, z84b2eb77e, z60a67f27d, zc44f0ab3b, ze64054cb6, z197a0495d)BEGIN CASE z197a0495d IS WHEN"000"=>pixd_out<=z163c5325c;WHEN"001"=>pixd_out<=z6bb6c7052;WHEN"010"=>pixd_out<=z0a9315da3;WHEN"011"=>pixd_out<=z564ee05a3;WHEN"100"=>pixd_out<=z84b2eb77e;WHEN"101"=>pixd_out<=z60a67f27d;WHEN"110"=>pixd_out<=zc44f0ab3b;WHEN"111"=>pixd_out<=ze64054cb6;WHEN OTHERS=>pixd_out<=(OTHERS=>'X');END CASE;END PROCESS z7d086e91c;zf5226fb5c<=y;z16921971f:PROCESS(zf5226fb5c)VARIABLE z925f2bf10:std_logic_vector(7 DOWNTO 0);BEGIN z925f2bf10:=zf5226fb5c(7 DOWNTO 0);z1934d98a3<=z925f2bf10(0);zb48298c48<=z925f2bf10(1);z75dc1577a<=z925f2bf10(2);z833ab3bd5<=z925f2bf10(3);z0068e7d64<=z925f2bf10(4);zb30429bb4<=z925f2bf10(5);z9f041aaff<=z925f2bf10(6);zcf058ee7c<=z925f2bf10(7);END PROCESS z16921971f;U_0:reg_bank_1px PORT MAP(clk=>clk,nullify=>nullify,pixd_in=>pixd_in,rst_n=>rst_n,write=>zc57c46db4,pixd_out=>z163c5325c);U_1:reg_bank_1px PORT MAP(clk=>clk,nullify=>nullify,pixd_in=>pixd_in,rst_n=>rst_n,write=>z1ea89dc0d,pixd_out=>z6bb6c7052);U_3:reg_bank_1px PORT MAP(clk=>clk,nullify=>nullify,pixd_in=>pixd_in,rst_n=>rst_n,write=>zcd48e1f4f,pixd_out=>z0a9315da3);U_4:reg_bank_1px PORT MAP(clk=>clk,nullify=>nullify,pixd_in=>pixd_in,rst_n=>rst_n,write=>z36424fa31,pixd_out=>z564ee05a3);U_5:reg_bank_1px PORT MAP(clk=>clk,nullify=>nullify,pixd_in=>pixd_in,rst_n=>rst_n,write=>z508ec0017,pixd_out=>z84b2eb77e);U_6:reg_bank_1px PORT MAP(clk=>clk,nullify=>nullify,pixd_in=>pixd_in,rst_n=>rst_n,write=>ze6d31b4ac,pixd_out=>z60a67f27d);U_11:reg_bank_1px PORT MAP(clk=>clk,nullify=>nullify,pixd_in=>pixd_in,rst_n=>rst_n,write=>z1b791bfd5,pixd_out=>zc44f0ab3b);U_12:reg_bank_1px PORT MAP(clk=>clk,nullify=>nullify,pixd_in=>pixd_in,rst_n=>rst_n,write=>z45a1dff88,pixd_out=>ze64054cb6);END struct;